// Created Tue Jan 20 16:49:41 2026

module nor_tb ();

  always begin

  end
endmodule
